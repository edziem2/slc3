module alu (
	input logic [15:0] A, B,
	input logic [1:0] ALUK,
	output logic [15:0] ALU_Out
);


endmodule 